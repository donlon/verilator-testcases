package mypkg;
    typedef int subtype_t;
endpackage
